--------------------------------------------------------------------------------
-- PROJECT: PIPE MANIA - GAME FOR FPGA
--------------------------------------------------------------------------------
-- NAME:    BRAM_ROM_SCREEN
-- AUTHORS: Tomáš Bannert <xbanne00@stud.feec.vutbr.cz>
-- LICENSE: The MIT License, please read LICENSE file
-- WEBSITE: https://github.com/jakubcabal/pipemania-fpga-game
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BRAM_ROM_SCREEN is
    Port (
        CLK      : in  std_logic;
        ROM_ADDR : in  std_logic_vector(11 downto 0);
        ROM_DOUT : out std_logic_vector(8 downto 0)
    );
end BRAM_ROM_SCREEN;

architecture FULL of BRAM_ROM_SCREEN is

    type rom_t is array (0 to 4095) of std_logic_vector(0 to 8);
    constant ROM : rom_t :=
    (
        -- main screen
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --1.r

        "000000000",
        "000000000",
        "000000000",
        "110010100",
        "000001100",
        "000010100",
        "000000000",
        "000011100",
        "000000000",
        "110010100",
        "000001100",
        "000010100",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --2.r

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --3.r

        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --4.r

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --5.r

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --6.r

        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --7.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --8.r

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --9.r

        "000011100",
        "000010100",
        "000000000",
        "110010100",
        "000011100",
        "000000000",
        "110010100",
        "000000000",
        "000010100",
        "000000000",
        "000011100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "110010100",
        "000000000",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --10.r

        "010001100",
        "000000000",
        "000001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "100010100",
        "000011100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --11.r

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000011100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000011100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --12.r

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --13.r

        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --14.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001001100",
        "001101100",
        "001110100",
        "001111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --15.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --16.r

        --game screen

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --1.r

        "000000000",
        "000110100",
        "000111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --2.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000101", -- KOMP0
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --3.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --4.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000110", -- KOMP1
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --5.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --6.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000111", -- KOMP2
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --7.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --8.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000001", -- KOMP3
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --9.r

        "000000000",
        "000101100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --10.r

        "000000000",
        "000100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000010", -- KOMP4
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --11.r

        "001011100",
        "001010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --12.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --13.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001000100",
        "000111100",
        "000111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --14.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --15.r

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --16.r
        -- win screen
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --1.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --2.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "110010100",
        "000001100",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --3.ř.

        "000000000",
        "000000000",
        "100010100",
        "000011100",
        "010010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --4.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "100010100",
        "000001100",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --5.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --6.ř.

        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --7.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --8.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "110010100",
        "000001100",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --9.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --10.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "100010100",
        "000011100",
        "000000000",
        "100010100",
        "000001100",
        "010010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --11.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --12.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "110010100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --13.ř.

        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "100010100",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --14.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --15.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000", --16.r
        -- lose screen
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --1.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --2.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "100010100",
        "010001100",
        "000010100",
        "110010100",
        "000001100",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --3.ř.

        "000000000",
        "000000000",
        "100010100",
        "000011100",
        "010010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "100010100",
        "000001100",
        "010010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --4.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "110010100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --5.ř.

        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "110010100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --6.ř.

        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "100010100",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --7.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --8.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000001100",
        "000001100",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --9.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --10.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --11.ř.

        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --12.ř.

        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000001100",
        "000000000",
        "000000000",
        "000001100",
        "000001100",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --13.ř.

        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --14.r.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --15.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --16.ř.
        -- lvl2
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --1.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --2.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --3.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --4.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --5.ř.

        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --6.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --7.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --8.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --9.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --10.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --11.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --12.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --13.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --14.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001001100",
        "001101100",
        "001110100",
        "001111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --15.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --16.ř.
        -- lvl3
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --1.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --2.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --3.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --4.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --5.ř.

        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --6.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --7.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --8.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --9.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --10.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --11.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --12.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --13.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --14.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001001100",
        "001101100",
        "001110100",
        "001111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --15.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --16.ř.
        -- lvl4
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --1.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000010100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --2.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --3.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "010001100",
        "000000000",
        "000011100",
        "000001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --4.ř.

        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --5.ř.

        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "010001100",
        "000000000",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000011100",
        "000001100",
        "010010100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --6.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --7.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --8.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --9.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --10.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --11.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --12.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --13.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001100100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --14.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "001001100",
        "001101100",
        "001110100",
        "001111100",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --15.ř.

        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",
        "000000000",   --16.ř.

        others => (others => '0')
    );

begin

    process (CLK)
    begin
        if (rising_edge(CLK)) then
            ROM_DOUT <= ROM(to_integer(unsigned(ROM_ADDR)));
        end if;
    end process;

end FULL;
