Z80_CMON_ROM_inst : Z80_CMON_ROM PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
