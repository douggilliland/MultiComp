---------------------------------------------------------------------------------------------
-- Taken from fpga4student.com
-- https://www.fpga4student.com/2017/09/vhdl-code-for-seven-segment-display.html
-- VHDL code for seven-segment display
-- Tested on A4-CE6 card
---------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
entity ElapsedTimeCounter_7S8D_LED  is
    Port ( clock_50Mhz : in STD_LOGIC;
           n_reset : in STD_LOGIC; -- active low reset
           Anode_Activate : out STD_LOGIC_VECTOR (7 downto 0);-- 8 Anode signals
           LED_out : out STD_LOGIC_VECTOR (7 downto 0));-- Cathode patterns of 7-segment display with Decimal Point
end ElapsedTimeCounter_7S8D_LED ;

architecture Behavioral of ElapsedTimeCounter_7S8D_LED  is
signal one_second_counter: STD_LOGIC_VECTOR (27 downto 0);
-- counter for generating 1-second clock enable
signal one_second_enable: std_logic;
-- one second enable for counting numbers
signal displayed_number: STD_LOGIC_VECTOR (31 downto 0);
-- counting decimal number to be displayed on 8-digit 7-segment display
signal LED_HEX: STD_LOGIC_VECTOR (3 downto 0);
signal refresh_counter: STD_LOGIC_VECTOR (20 downto 0);
-- creating 10.5ms refresh period
signal LED_activating_counter: std_logic_vector(2 downto 0);
-- the other 3-bit for creating 8 LED-activating signals
-- count         0		->  1  ->  2  ->  3 -> 4 -> 5 -> 6 -> 7
-- activates    LED1	LED2   LED3   LED4
-- and repeat
begin
-- VHDL code for Hex to 7-segment decoder
-- Cathode patterns of the 7-segment LED display 
process(LED_HEX)
begin
    case LED_HEX is
    when x"0" => LED_out <= "11000000"; -- "0" - bit order is dp - g thru a
    when x"1" => LED_out <= "11111001"; -- "1" 
    when x"2" => LED_out <= "10100100"; -- "2" 
    when x"3" => LED_out <= "10110000"; -- "3" 
    when x"4" => LED_out <= "10011001"; -- "4" 
    when x"5" => LED_out <= "10010010"; -- "5" 
    when x"6" => LED_out <= "10000010"; -- "6" 
    when x"7" => LED_out <= "11111000"; -- "7" 
    when x"8" => LED_out <= "10000000"; -- "8"     
    when x"9" => LED_out <= "10010000"; -- "9" 
    when x"A" => LED_out <= "10001000"; -- "A"
    when x"B" => LED_out <= "10000011"; -- "B"
    when x"C" => LED_out <= "11000110"; -- "C"
    when x"D" => LED_out <= "10100001"; -- "D"
    when x"E" => LED_out <= "10000110"; -- "E"
    when x"F" => LED_out <= "10001110"; -- "F"
    end case;
end process;
-- 7-segment display controller
-- generate refresh period of 10.5ms
process(clock_50Mhz,n_reset)
begin 
    if(n_reset='0') then
        refresh_counter <= (others => '0');
    elsif(rising_edge(clock_50Mhz)) then
        refresh_counter <= refresh_counter + 1;
    end if;
end process;
 LED_activating_counter <= refresh_counter(19 downto 17);
-- 4-to-1 MUX to generate anode activating signals for 4 LEDs 
process(LED_activating_counter)
begin
    case LED_activating_counter is
    when "000" =>
        Anode_Activate <= "11111110"; 
        -- activate LED1 and Deactivate LED2, LED3, LED4
        LED_HEX <= displayed_number(31 downto 28);
        -- the first hex digit of the 16-bit number
    when "001" =>
        Anode_Activate <= "11111101"; 
        -- activate LED2 and Deactivate LED1, LED3, LED4
        LED_HEX <= displayed_number(27 downto 24);
        -- the second hex digit of the 16-bit number
    when "010" =>
        Anode_Activate <= "11111011"; 
        -- activate LED3 and Deactivate LED2, LED1, LED4
        LED_HEX <= displayed_number(23 downto 20);
        -- the third hex digit of the 16-bit number
    when "011" =>
        Anode_Activate <= "11110111"; 
        -- activate LED4 and Deactivate LED2, LED3, LED1
        LED_HEX <= displayed_number(19 downto 16);
        -- the fourth hex digit of the 16-bit number    
    when "100" =>
        Anode_Activate <= "11101111"; 
        -- activate LED5 and Deactivate LED2, LED3, LED4
        LED_HEX <= displayed_number(15 downto 12);
        -- the first hex digit of the 16-bit number
    when "101" =>
        Anode_Activate <= "11011111"; 
        -- activate LED6 and Deactivate LED1, LED3, LED4
        LED_HEX <= displayed_number(11 downto 8);
        -- the second hex digit of the 16-bit number
    when "110" =>
        Anode_Activate <= "10111111"; 
        -- activate LED7 and Deactivate LED2, LED1, LED4
        LED_HEX <= displayed_number(7 downto 4);
        -- the third hex digit of the 16-bit number
    when "111" =>
        Anode_Activate <= "01111111"; 
        -- activate LED8 and Deactivate LED2, LED3, LED1
        LED_HEX <= displayed_number(3 downto 0);
        -- the fourth hex digit of the 16-bit number    
    end case;
end process;
-- Counting the number to be displayed on 8-digit 7-segment Display 
-- on Basys 3 FPGA board
process(clock_50Mhz, n_reset)
begin
        if(n_reset='0') then
            one_second_counter <= (others => '0');
        elsif(rising_edge(clock_50Mhz)) then
            if(one_second_counter>=x"2FAF07F") then
                one_second_counter <= (others => '0');
            else
                one_second_counter <= one_second_counter + "0000001";
            end if;
        end if;
end process;
one_second_enable <= '1' when one_second_counter=x"2FAF07F" else '0';
process(clock_50Mhz, n_reset)
begin
        if(n_reset='0') then
            displayed_number <= (others => '0');
        elsif(rising_edge(clock_50Mhz)) then
             if(one_second_enable='1') then
                displayed_number <= displayed_number + x"00000001";
             end if;
        end if;
end process;
end Behavioral;
