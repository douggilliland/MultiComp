library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY CharRom IS
	PORT
	(
		address : in std_logic_vector(10 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END CharRom;

architecture behavior of CharRom is
type romtable is array (0 to 2047) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"5A",x"7E",x"5A",x"18",x"18",x"5A",x"7E",x"5A",x"42",x"7E",x"5A",x"18",x"18",x"5A",x"7E",x"42",x"81",x"42",x"24",x"24",x"24",x"24",x"42",x"81",x"81",x"42",x"3C",x"00",x"00",x"3C",x"42",x"81",
x"00",x"00",x"00",x"24",x"99",x"5A",x"FF",x"00",x"FF",x"FF",x"C3",x"C3",x"00",x"00",x"00",x"00",x"FF",x"FF",x"C3",x"C3",x"C3",x"C3",x"FF",x"FF",x"00",x"00",x"00",x"00",x"C3",x"C3",x"FF",x"FF",
x"FF",x"FF",x"C3",x"DB",x"DB",x"C3",x"FF",x"FF",x"18",x"24",x"24",x"42",x"42",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"28",x"44",x"00",x"00",x"00",
x"00",x"00",x"F8",x"00",x"F8",x"00",x"F8",x"00",x"18",x"3C",x"7E",x"7F",x"7E",x"3C",x"08",x"08",x"00",x"00",x"18",x"3C",x"7E",x"7E",x"56",x"5E",x"18",x"3D",x"7F",x"FF",x"AD",x"FF",x"AD",x"BF",
x"18",x"3C",x"5A",x"18",x"18",x"18",x"18",x"3C",x"0F",x"07",x"0F",x"1D",x"B8",x"70",x"20",x"10",x"00",x"04",x"82",x"FF",x"FF",x"82",x"04",x"00",x"10",x"20",x"70",x"B8",x"1D",x"0F",x"07",x"0F",
x"3C",x"18",x"18",x"18",x"18",x"5A",x"3C",x"18",x"08",x"04",x"0E",x"1D",x"B8",x"F0",x"E0",x"F0",x"00",x"20",x"41",x"FF",x"FF",x"41",x"20",x"00",x"F0",x"E0",x"F0",x"B8",x"1D",x"0E",x"04",x"08",
x"18",x"24",x"20",x"70",x"20",x"20",x"7C",x"00",x"00",x"00",x"00",x"02",x"7E",x"40",x"00",x"00",x"00",x"38",x"28",x"28",x"7C",x"28",x"38",x"00",x"00",x"38",x"28",x"28",x"28",x"28",x"38",x"00",
x"10",x"70",x"F0",x"70",x"10",x"00",x"00",x"00",x"18",x"24",x"42",x"81",x"18",x"24",x"42",x"81",x"00",x"7E",x"42",x"24",x"18",x"18",x"18",x"18",x"81",x"42",x"24",x"18",x"81",x"42",x"24",x"18",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"00",x"28",x"28",x"28",x"00",x"00",x"00",x"00",x"00",x"28",x"28",x"7C",x"28",x"7C",x"28",x"28",x"00",
x"10",x"3C",x"50",x"38",x"14",x"78",x"10",x"00",x"60",x"64",x"08",x"10",x"20",x"4C",x"0C",x"00",x"20",x"50",x"50",x"20",x"54",x"48",x"34",x"00",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",
x"10",x"20",x"40",x"40",x"40",x"20",x"10",x"00",x"10",x"08",x"04",x"04",x"04",x"08",x"10",x"00",x"10",x"54",x"38",x"10",x"38",x"54",x"10",x"00",x"00",x"10",x"10",x"7C",x"10",x"10",x"00",x"00",
x"00",x"00",x"00",x"00",x"10",x"10",x"20",x"00",x"00",x"00",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"00",x"04",x"08",x"10",x"20",x"40",x"00",x"00",
x"38",x"44",x"4C",x"54",x"64",x"44",x"38",x"00",x"10",x"30",x"10",x"10",x"10",x"10",x"38",x"00",x"38",x"44",x"04",x"18",x"20",x"40",x"7C",x"00",x"7C",x"04",x"08",x"18",x"04",x"44",x"38",x"00",
x"08",x"18",x"28",x"48",x"7C",x"08",x"08",x"00",x"7C",x"40",x"78",x"04",x"04",x"44",x"38",x"00",x"1C",x"20",x"40",x"78",x"44",x"44",x"38",x"00",x"7C",x"04",x"08",x"10",x"20",x"20",x"20",x"00",
x"38",x"44",x"44",x"38",x"44",x"44",x"38",x"00",x"38",x"44",x"44",x"3C",x"04",x"08",x"70",x"00",x"00",x"00",x"10",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"10",x"10",x"20",x"00",
x"08",x"10",x"20",x"40",x"20",x"10",x"08",x"00",x"00",x"00",x"7C",x"00",x"7C",x"00",x"00",x"00",x"20",x"10",x"08",x"04",x"08",x"10",x"20",x"00",x"38",x"44",x"08",x"10",x"10",x"00",x"10",x"00",
x"38",x"44",x"54",x"5C",x"58",x"40",x"3C",x"00",x"10",x"28",x"44",x"44",x"7C",x"44",x"44",x"00",x"78",x"44",x"44",x"78",x"44",x"44",x"78",x"00",x"38",x"44",x"40",x"40",x"40",x"44",x"38",x"00",
x"78",x"44",x"44",x"44",x"44",x"44",x"78",x"00",x"7C",x"40",x"40",x"78",x"40",x"40",x"7C",x"00",x"7C",x"40",x"40",x"78",x"40",x"40",x"40",x"00",x"3C",x"40",x"40",x"40",x"4C",x"44",x"3C",x"00",
x"44",x"44",x"44",x"7C",x"44",x"44",x"44",x"00",x"38",x"10",x"10",x"10",x"10",x"10",x"38",x"00",x"04",x"04",x"04",x"04",x"04",x"44",x"38",x"00",x"44",x"48",x"50",x"60",x"50",x"48",x"44",x"00",
x"40",x"40",x"40",x"40",x"40",x"40",x"7C",x"00",x"44",x"6C",x"54",x"54",x"44",x"44",x"44",x"00",x"44",x"44",x"64",x"54",x"4C",x"44",x"44",x"00",x"38",x"44",x"44",x"44",x"44",x"44",x"38",x"00",
x"78",x"44",x"44",x"78",x"40",x"40",x"40",x"00",x"38",x"44",x"44",x"44",x"54",x"48",x"34",x"00",x"78",x"44",x"44",x"78",x"50",x"48",x"44",x"00",x"38",x"44",x"40",x"38",x"04",x"44",x"38",x"00",
x"7C",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"38",x"00",x"44",x"44",x"44",x"44",x"44",x"28",x"10",x"00",x"44",x"44",x"44",x"54",x"54",x"6C",x"44",x"00",
x"44",x"44",x"28",x"10",x"28",x"44",x"44",x"00",x"44",x"44",x"28",x"10",x"10",x"10",x"10",x"00",x"7C",x"04",x"08",x"10",x"20",x"40",x"7C",x"00",x"7C",x"60",x"60",x"60",x"60",x"60",x"7C",x"00",
x"00",x"40",x"20",x"10",x"08",x"04",x"00",x"00",x"7C",x"0C",x"0C",x"0C",x"0C",x"0C",x"7C",x"00",x"10",x"38",x"54",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"34",x"4C",x"44",x"4C",x"34",x"00",x"40",x"40",x"58",x"64",x"44",x"64",x"58",x"00",x"00",x"00",x"3C",x"40",x"40",x"40",x"3C",x"00",
x"04",x"04",x"34",x"4C",x"44",x"4C",x"34",x"00",x"00",x"00",x"38",x"44",x"7C",x"40",x"38",x"00",x"08",x"10",x"10",x"38",x"10",x"10",x"10",x"00",x"00",x"34",x"4C",x"44",x"4C",x"34",x"04",x"38",
x"40",x"40",x"78",x"44",x"44",x"44",x"44",x"00",x"00",x"10",x"00",x"30",x"10",x"10",x"38",x"00",x"00",x"08",x"00",x"08",x"08",x"08",x"08",x"30",x"40",x"44",x"48",x"50",x"70",x"48",x"44",x"00",
x"30",x"10",x"10",x"10",x"10",x"10",x"38",x"00",x"00",x"00",x"68",x"54",x"54",x"54",x"54",x"00",x"00",x"00",x"78",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"38",x"44",x"44",x"44",x"38",x"00",
x"00",x"58",x"64",x"44",x"64",x"58",x"40",x"40",x"00",x"34",x"4C",x"44",x"4C",x"34",x"04",x"04",x"00",x"00",x"58",x"60",x"40",x"40",x"40",x"00",x"00",x"00",x"3C",x"40",x"38",x"04",x"78",x"00",
x"00",x"10",x"7C",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"3C",x"00",x"00",x"00",x"44",x"44",x"28",x"28",x"10",x"00",x"00",x"00",x"44",x"44",x"44",x"54",x"28",x"00",
x"00",x"00",x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"00",x"24",x"24",x"24",x"3C",x"04",x"38",x"00",x"00",x"7C",x"08",x"10",x"20",x"7C",x"00",x"0C",x"10",x"10",x"20",x"10",x"10",x"0C",x"00",
x"60",x"10",x"10",x"08",x"10",x"10",x"60",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"00",x"00",x"10",x"00",x"7C",x"00",x"10",x"00",x"00",x"00",x"00",x"04",x"38",x"40",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",
x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",
x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",
x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"00",x"10",x"08",x"FC",x"02",x"FC",x"08",x"10",
x"00",x"10",x"20",x"7E",x"80",x"7E",x"20",x"10",x"00",x"00",x"28",x"7C",x"82",x"7C",x"28",x"00",x"00",x"00",x"10",x"28",x"44",x"FE",x"00",x"00",x"AA",x"55",x"AA",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"AA",x"55",x"AA",x"55",x"A0",x"50",x"A0",x"50",x"A0",x"50",x"A0",x"50",x"0A",x"05",x"0A",x"05",x"0A",x"05",x"0A",x"05",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",
x"81",x"42",x"24",x"18",x"18",x"24",x"42",x"81",x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"81",x"42",x"24",x"18",x"00",x"00",x"00",x"00",
x"01",x"02",x"04",x"08",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"00",x"18",x"24",x"42",x"81",x"80",x"40",x"20",x"10",x"10",x"20",x"40",x"80",x"03",x"0C",x"30",x"C0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"03",x"0C",x"30",x"C0",x"C0",x"30",x"0C",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"30",x"0C",x"03",x"08",x"08",x"04",x"04",x"02",x"02",x"01",x"01",
x"80",x"80",x"40",x"40",x"20",x"20",x"10",x"10",x"01",x"01",x"02",x"02",x"04",x"04",x"08",x"08",x"10",x"10",x"20",x"20",x"40",x"40",x"80",x"80",x"08",x"08",x"08",x"0F",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"0F",x"08",x"08",x"08",x"00",x"00",x"00",x"00",x"F0",x"10",x"10",x"10",x"10",x"10",x"10",x"F0",x"00",x"00",x"00",x"00",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"1C",x"10",x"10",x"10",x"50",x"30",x"10",x"00",
x"08",x"14",x"10",x"10",x"10",x"50",x"20",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"10",x"2A",x"04",x"10",x"2A",x"04",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",
x"18",x"18",x"18",x"1F",x"1F",x"18",x"18",x"18",x"00",x"00",x"00",x"FF",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"F8",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",
x"08",x"08",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"04",x"08",x"08",x"00",x"00",x"00",x"00",x"C0",x"20",x"10",x"10",x"10",x"10",x"20",x"C0",x"00",x"00",x"00",x"00",
x"03",x"04",x"08",x"08",x"08",x"08",x"04",x"03",x"C0",x"20",x"10",x"10",x"10",x"10",x"20",x"C0",x"3C",x"42",x"81",x"81",x"81",x"81",x"42",x"3C",x"0F",x"30",x"C0",x"C0",x"C0",x"C0",x"30",x"0F",
x"F0",x"0C",x"03",x"03",x"03",x"03",x"0C",x"F0",x"00",x"66",x"FF",x"FF",x"7E",x"3C",x"18",x"00",x"1C",x"1C",x"6B",x"7F",x"6B",x"08",x"08",x"08",x"18",x"3C",x"7E",x"FF",x"FF",x"18",x"18",x"3C",
x"18",x"3C",x"7E",x"FF",x"7E",x"3C",x"18",x"00",x"E7",x"C3",x"81",x"00",x"00",x"81",x"C3",x"E7",x"03",x"0F",x"3F",x"FF",x"FF",x"3F",x"0F",x"03",x"C0",x"F0",x"FC",x"FF",x"FF",x"FC",x"F0",x"C0",
x"18",x"18",x"3C",x"7E",x"FF",x"DB",x"18",x"3C",x"30",x"38",x"9C",x"FF",x"FF",x"9C",x"38",x"30",x"3C",x"18",x"DB",x"FF",x"7E",x"3C",x"18",x"18",x"0C",x"1C",x"39",x"FF",x"FF",x"39",x"1C",x"0C",
x"00",x"00",x"00",x"10",x"38",x"54",x"10",x"28",x"00",x"00",x"00",x"34",x"48",x"48",x"34",x"00",x"18",x"24",x"24",x"38",x"24",x"24",x"38",x"40",x"00",x"00",x"00",x"28",x"44",x"54",x"28",x"00",
x"38",x"40",x"40",x"30",x"48",x"48",x"30",x"00",x"10",x"10",x"54",x"54",x"38",x"10",x"10",x"00",x"00",x"00",x"38",x"44",x"44",x"28",x"C6",x"00",x"00",x"24",x"24",x"24",x"38",x"20",x"20",x"00",
x"00",x"00",x"3C",x"68",x"28",x"28",x"28",x"00",x"7C",x"20",x"10",x"18",x"10",x"20",x"7C",x"00",x"00",x"00",x"40",x"20",x"10",x"28",x"44",x"00",x"10",x"10",x"38",x"54",x"54",x"38",x"10",x"00",
x"38",x"44",x"44",x"7C",x"44",x"44",x"38",x"00",x"00",x"00",x"18",x"20",x"38",x"20",x"18",x"00",x"00",x"00",x"64",x"24",x"28",x"30",x"20",x"00",x"00",x"00",x"64",x"18",x"10",x"30",x"30",x"00"
);
begin
process (address)
begin
q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;

