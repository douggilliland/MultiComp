--------------------------------------------------------------------------------
-- PROJECT: PIPE MANIA - GAME FOR FPGA
--------------------------------------------------------------------------------
-- NAME:    BRAM_ROM_CELL
-- AUTHORS: Tomáš Bannert <xbanne00@stud.feec.vutbr.cz>
-- LICENSE: The MIT License, please read LICENSE file
-- WEBSITE: https://github.com/jakubcabal/pipemania-fpga-game
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BRAM_ROM_CELL is
    Port (
        CLK      : in  std_logic;
        ROM_ADDR : in  std_logic_vector(8 downto 0);
        ROM_DOUT : out std_logic_vector(31 downto 0)
    );
end BRAM_ROM_CELL;

architecture FULL of BRAM_ROM_CELL is

    type rom_t is array (0 to 511) of std_logic_vector(0 to 31);
    constant ROM : rom_t :=
    (
        "11111111111111111111111111111111",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "10000000000000000000000000000001",
        "11111111111111111111111111111111",

        -- Dalsi obrazek (rovna 1=modra) -- 0001

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- Dalsi obrazek (zahnuta 1=modra) 0010

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11100000000000000000000000000000",
        "11100000000000000000000000000000",
        "11100000000000000000000000000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "11111111111111111111111110000000",
        "00000000000000001111111110000000",
        "00000000000000001111111110000000",
        "00000000000000000011111110000000",
        "00000000000000000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11111111111111000011111110000000",
        "11100001111111000011111110000000",
        "11100001111111000011111110000000",
        "11100001111111000011111110000000",
        "00000001111111000011111110000000",
        "00001111111111000011111111110000",
        "00001111111111000011111111110000",
        "00001111111111000011111111110000",

        -- Dalsi obrazek (T 1=modra) - 0011

        "00001111111111000011111111110000",
        "00001111111111000011111111110000",
        "00001111111111000011111111110000",
        "00000001111111000011111110000000",
        "11100001111111000011111110000111",
        "11100001111111000011111110000111",
        "11100001111111000011111110000111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11111111111111000011111111111111",
        "11100001111111000011111110000111",
        "11100001111111000011111110000111",
        "11100001111111000011111110000111",
        "00000001111111000011111110000000",
        "00001111111111000011111111110000",
        "00001111111111000011111111110000",
        "00001111111111000011111111110000",

        -- Dalsi obrazek (spodni cast bocni trubky 1=modra) - 0100

        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111001110011100111001110011111",
        "11111001110011100111001110011111",
        "01111111111111111111111111111110",
        "01111111111111111111111111111110",
        "01111111111111111111111111111110",
        "00111111111111111111111111111100",
        "00111111111111111111111111111100",
        "00011111111111111111111111111000",
        "00001111111111111111111111110000",
        "00000111111111111111111111100000",
        "00000011111111111111111111000000",
        "00000001111111111111111110000000",
        "00000000011111111111111000000000",
        "00000000000011111111000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",

        -- Dalsi obrazek (telo trubky 1=bila 8x) - 0101

        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",
        "00100000000000000000000000000100",


        -- Dalsi obrazek (vrchni cast bocni trubky 1=modra) - 0110

        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",

        -- Dalsi obrazek (propojka bocni trubky s hernim polem 1=modra) - 0111

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- Dalsi obrazek (koncova trubka 1=modra) - 1000

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111000011111111111111",
        "11111111111100111100111111111111",
        "11111111111001111110011111111111",
        "11111111111010111101011111111111",
        "11111111110111011011101111111111",
        "11111111110111100111101111111111",
        "11111111110111100111101111111111",
        "11111111110111011011101111111111",
        "11111111111010111101011111111111",
        "11111111111001111110011111111111",
        "11111111111100111100111111111111",
        "11111111111111000011111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11100000000000000000000000000111",
        "11100000000000000000000000000111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- text1 (bila) - 1001

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00011110000111100001111110000111",
        "00011110000111100001111110000111",
        "00011001100110011001100000011000",
        "00011001100110011001100000011000",
        "00011110000111100001111000000110",
        "00011110000111100001111000000110",
        "00011000000110011001100000000001",
        "00011000000110011001100000000001",
        "00011000000110011001111110011110",
        "00011000000110011001111110011110",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000001100001",
        "00000000000000000000000001100001",
        "00000000000000000000000110011001",
        "00000000000000000000000110011001",
        "00000000000000000000000110011001",
        "00000000000000000000000110011001",
        "00000000000000000000000110011001",
        "00000000000000000000000110011001",
        "00000000000000000000000001100001",
        "00000000000000000000000001100001",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- Dalsi obrazek (tenka trubka ke startovni ohnuta 1=modra) - 1010

        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000",
        "00000000000001111100000000000000",
        "00000000000011111100000000000000",
        "11111111111111111000000000000000",
        "11111111111111111000000000000000",
        "11111111111111110000000000000000",
        "11111111111111000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- Dalsi obrazek (tenka trubka ke startovni rovna 1=modra) - 1011

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- Dalsi obrazek (cihla 1=cervena) - 1100

        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "00000000000000000000000000000000",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "00000000000000000000000000000000",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "00000000000000000000000000000000",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "00000000000000000000000000000000",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "00000000000000000000000000000000",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "00000000000000000000000000000000",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "01111111011111110111111101111111",
        "00000000000000000000000000000000",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "11110111111101111111011111110111",
        "00000000000000000000000000000000",

        -- text2 (bila) - 1101

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000011000000000011000",
        "00000000000000011000000000011000",
        "10000111100000011000011110011000",
        "10000111100000011000011110011000",
        "00011000000000000001100000000000",
        "00011000000000000001100000000000",
        "00000110000000000000011000000000",
        "00000110000000000000011000000000",
        "10000001100000000000000110000000",
        "10000001100000000000000110000000",
        "00011110000000000001111000000000",
        "00011110000000000001111000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11100001100110011000011000011001",
        "11100001100110011000011000011001",
        "10011001100110011001100110011001",
        "10011001100110011001100110011001",
        "11100001100110011001100110011001",
        "11100001100110011001100110011001",
        "10011000011000011001100110011001",
        "10011000011000011001100110011001",
        "11100000011000011000011000000110",
        "11100000011000011000011000000110",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- text3 (bila) - 1110

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00011111100001100000000001111001",
        "00011111100001100000000001111001",
        "00000110000110011000000110000000",
        "00000110000110011000000110000000",
        "00000110000110011000000001100000",
        "00000110000110011000000001100000",
        "00000110000110011000000000011000",
        "00000110000110011000000000011000",
        "00000110000001100000000111100000",
        "00000110000001100000000111100000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000111100110000001100110000000",
        "00000111100110000001100110000000",
        "00011000000110000001100110000000",
        "00011000000110000001100110000000",
        "00000110000110000000011000000000",
        "00000110000110000000011000000000",
        "00000001100110000000011000000000",
        "00000001100110000000011000000000",
        "00011110000111111000011000011000",
        "00011110000111111000011000011000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        -- text4 (bila) - 1111

        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "11111000011000011110000111111000",
        "11111000011000011110000111111000",
        "01100001100110011001100001100000",
        "01100001100110011001100001100000",
        "01100001100110011110000001100000",
        "01100001100110011110000001100000",
        "01100001111110011001100001100000",
        "01100001111110011001100001100000",
        "01100001100110011001100001100000",
        "01100001100110011001100001100000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00011000000000000000000000000000",
        "00011000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",

        others => (others => '0')
    );

begin

    process (CLK)
    begin
        if (rising_edge(CLK)) then
            ROM_DOUT <= ROM(to_integer(unsigned(ROM_ADDR)));
        end if;
    end process;

end FULL;
